// nios.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module nios (
		output wire       arbitrotx_writeresponsevalid_n,           //                      arbitrotx.writeresponsevalid_n
		input  wire       clk_clk,                                  //                            clk.clk
		output wire [7:0] lcd_0_conduit_end_1_readdata,             //            lcd_0_conduit_end_1.readdata
		output wire       lcd_0_conduit_end_2_writeresponsevalid_n, //            lcd_0_conduit_end_2.writeresponsevalid_n
		output wire       lcd_0_conduit_end_3_writeresponsevalid_n, //            lcd_0_conduit_end_3.writeresponsevalid_n
		output wire       lcd_0_conduit_end_4_writeresponsevalid_n, //            lcd_0_conduit_end_4.writeresponsevalid_n
		output wire [3:0] leds_external_connection_export,          //       leds_external_connection.export
		input  wire [3:0] pushbutton_external_connection_export,    // pushbutton_external_connection.export
		input  wire       uart_0_external_connection_rxd,           //     uart_0_external_connection.rxd
		output wire       uart_0_external_connection_txd            //                               .txd
	);

	wire         nios2_debug_reset_request_reset;                                          // nios2:debug_reset_request -> [rst_controller:reset_in0, rst_controller:reset_in1]
	wire         nios2_custom_instruction_master_readra;                                   // nios2:D_ci_readra -> nios2_custom_instruction_master_translator:ci_slave_readra
	wire   [4:0] nios2_custom_instruction_master_a;                                        // nios2:D_ci_a -> nios2_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] nios2_custom_instruction_master_b;                                        // nios2:D_ci_b -> nios2_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] nios2_custom_instruction_master_c;                                        // nios2:D_ci_c -> nios2_custom_instruction_master_translator:ci_slave_c
	wire         nios2_custom_instruction_master_readrb;                                   // nios2:D_ci_readrb -> nios2_custom_instruction_master_translator:ci_slave_readrb
	wire         nios2_custom_instruction_master_clk;                                      // nios2:E_ci_multi_clock -> nios2_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] nios2_custom_instruction_master_ipending;                                 // nios2:W_ci_ipending -> nios2_custom_instruction_master_translator:ci_slave_ipending
	wire         nios2_custom_instruction_master_start;                                    // nios2:E_ci_multi_start -> nios2_custom_instruction_master_translator:ci_slave_multi_start
	wire         nios2_custom_instruction_master_reset_req;                                // nios2:E_ci_multi_reset_req -> nios2_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios2_custom_instruction_master_done;                                     // nios2_custom_instruction_master_translator:ci_slave_multi_done -> nios2:E_ci_multi_done
	wire   [7:0] nios2_custom_instruction_master_n;                                        // nios2:D_ci_n -> nios2_custom_instruction_master_translator:ci_slave_n
	wire  [31:0] nios2_custom_instruction_master_result;                                   // nios2_custom_instruction_master_translator:ci_slave_result -> nios2:E_ci_result
	wire         nios2_custom_instruction_master_estatus;                                  // nios2:W_ci_estatus -> nios2_custom_instruction_master_translator:ci_slave_estatus
	wire         nios2_custom_instruction_master_clk_en;                                   // nios2:E_ci_multi_clk_en -> nios2_custom_instruction_master_translator:ci_slave_multi_clken
	wire  [31:0] nios2_custom_instruction_master_datab;                                    // nios2:E_ci_datab -> nios2_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] nios2_custom_instruction_master_dataa;                                    // nios2:E_ci_dataa -> nios2_custom_instruction_master_translator:ci_slave_dataa
	wire         nios2_custom_instruction_master_reset;                                    // nios2:E_ci_multi_reset -> nios2_custom_instruction_master_translator:ci_slave_multi_reset
	wire         nios2_custom_instruction_master_writerc;                                  // nios2:D_ci_writerc -> nios2_custom_instruction_master_translator:ci_slave_writerc
	wire         nios2_custom_instruction_master_translator_multi_ci_master_readra;        // nios2_custom_instruction_master_translator:multi_ci_master_readra -> nios2_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] nios2_custom_instruction_master_translator_multi_ci_master_a;             // nios2_custom_instruction_master_translator:multi_ci_master_a -> nios2_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] nios2_custom_instruction_master_translator_multi_ci_master_b;             // nios2_custom_instruction_master_translator:multi_ci_master_b -> nios2_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         nios2_custom_instruction_master_translator_multi_ci_master_clk;           // nios2_custom_instruction_master_translator:multi_ci_master_clk -> nios2_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios2_custom_instruction_master_translator_multi_ci_master_readrb;        // nios2_custom_instruction_master_translator:multi_ci_master_readrb -> nios2_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] nios2_custom_instruction_master_translator_multi_ci_master_c;             // nios2_custom_instruction_master_translator:multi_ci_master_c -> nios2_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         nios2_custom_instruction_master_translator_multi_ci_master_start;         // nios2_custom_instruction_master_translator:multi_ci_master_start -> nios2_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         nios2_custom_instruction_master_translator_multi_ci_master_reset_req;     // nios2_custom_instruction_master_translator:multi_ci_master_reset_req -> nios2_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios2_custom_instruction_master_translator_multi_ci_master_done;          // nios2_custom_instruction_master_multi_xconnect:ci_slave_done -> nios2_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios2_custom_instruction_master_translator_multi_ci_master_n;             // nios2_custom_instruction_master_translator:multi_ci_master_n -> nios2_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] nios2_custom_instruction_master_translator_multi_ci_master_result;        // nios2_custom_instruction_master_multi_xconnect:ci_slave_result -> nios2_custom_instruction_master_translator:multi_ci_master_result
	wire         nios2_custom_instruction_master_translator_multi_ci_master_clk_en;        // nios2_custom_instruction_master_translator:multi_ci_master_clken -> nios2_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] nios2_custom_instruction_master_translator_multi_ci_master_datab;         // nios2_custom_instruction_master_translator:multi_ci_master_datab -> nios2_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] nios2_custom_instruction_master_translator_multi_ci_master_dataa;         // nios2_custom_instruction_master_translator:multi_ci_master_dataa -> nios2_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios2_custom_instruction_master_translator_multi_ci_master_reset;         // nios2_custom_instruction_master_translator:multi_ci_master_reset -> nios2_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         nios2_custom_instruction_master_translator_multi_ci_master_writerc;       // nios2_custom_instruction_master_translator:multi_ci_master_writerc -> nios2_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_readra;         // nios2_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_a;              // nios2_custom_instruction_master_multi_xconnect:ci_master0_a -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_b;              // nios2_custom_instruction_master_multi_xconnect:ci_master0_b -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb;         // nios2_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_c;              // nios2_custom_instruction_master_multi_xconnect:ci_master0_c -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_clk;            // nios2_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending;       // nios2_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_start;          // nios2_custom_instruction_master_multi_xconnect:ci_master0_start -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req;      // nios2_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_done;           // nios2_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios2_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_n;              // nios2_custom_instruction_master_multi_xconnect:ci_master0_n -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_result;         // nios2_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios2_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus;        // nios2_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en;         // nios2_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_datab;          // nios2_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa;          // nios2_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_reset;          // nios2_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc;        // nios2_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk;    // nios2_custom_instruction_master_multi_slave_translator0:ci_master_clk -> LCD_0:clk
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en; // nios2_custom_instruction_master_multi_slave_translator0:ci_master_clken -> LCD_0:clk_en
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab;  // nios2_custom_instruction_master_multi_slave_translator0:ci_master_datab -> LCD_0:datab
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa;  // nios2_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> LCD_0:dataa
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_readra;         // nios2_custom_instruction_master_multi_xconnect:ci_master1_readra -> nios2_custom_instruction_master_multi_slave_translator1:ci_slave_readra
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master1_a;              // nios2_custom_instruction_master_multi_xconnect:ci_master1_a -> nios2_custom_instruction_master_multi_slave_translator1:ci_slave_a
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master1_b;              // nios2_custom_instruction_master_multi_xconnect:ci_master1_b -> nios2_custom_instruction_master_multi_slave_translator1:ci_slave_b
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_readrb;         // nios2_custom_instruction_master_multi_xconnect:ci_master1_readrb -> nios2_custom_instruction_master_multi_slave_translator1:ci_slave_readrb
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master1_c;              // nios2_custom_instruction_master_multi_xconnect:ci_master1_c -> nios2_custom_instruction_master_multi_slave_translator1:ci_slave_c
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_clk;            // nios2_custom_instruction_master_multi_xconnect:ci_master1_clk -> nios2_custom_instruction_master_multi_slave_translator1:ci_slave_clk
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master1_ipending;       // nios2_custom_instruction_master_multi_xconnect:ci_master1_ipending -> nios2_custom_instruction_master_multi_slave_translator1:ci_slave_ipending
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_start;          // nios2_custom_instruction_master_multi_xconnect:ci_master1_start -> nios2_custom_instruction_master_multi_slave_translator1:ci_slave_start
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_reset_req;      // nios2_custom_instruction_master_multi_xconnect:ci_master1_reset_req -> nios2_custom_instruction_master_multi_slave_translator1:ci_slave_reset_req
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_done;           // nios2_custom_instruction_master_multi_slave_translator1:ci_slave_done -> nios2_custom_instruction_master_multi_xconnect:ci_master1_done
	wire   [7:0] nios2_custom_instruction_master_multi_xconnect_ci_master1_n;              // nios2_custom_instruction_master_multi_xconnect:ci_master1_n -> nios2_custom_instruction_master_multi_slave_translator1:ci_slave_n
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master1_result;         // nios2_custom_instruction_master_multi_slave_translator1:ci_slave_result -> nios2_custom_instruction_master_multi_xconnect:ci_master1_result
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_estatus;        // nios2_custom_instruction_master_multi_xconnect:ci_master1_estatus -> nios2_custom_instruction_master_multi_slave_translator1:ci_slave_estatus
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_clk_en;         // nios2_custom_instruction_master_multi_xconnect:ci_master1_clken -> nios2_custom_instruction_master_multi_slave_translator1:ci_slave_clken
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master1_datab;          // nios2_custom_instruction_master_multi_xconnect:ci_master1_datab -> nios2_custom_instruction_master_multi_slave_translator1:ci_slave_datab
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master1_dataa;          // nios2_custom_instruction_master_multi_xconnect:ci_master1_dataa -> nios2_custom_instruction_master_multi_slave_translator1:ci_slave_dataa
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_reset;          // nios2_custom_instruction_master_multi_xconnect:ci_master1_reset -> nios2_custom_instruction_master_multi_slave_translator1:ci_slave_reset
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_writerc;        // nios2_custom_instruction_master_multi_xconnect:ci_master1_writerc -> nios2_custom_instruction_master_multi_slave_translator1:ci_slave_writerc
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator1_ci_master_result; // arbitro_0:result -> nios2_custom_instruction_master_multi_slave_translator1:ci_master_result
	wire         nios2_custom_instruction_master_multi_slave_translator1_ci_master_clk;    // nios2_custom_instruction_master_multi_slave_translator1:ci_master_clk -> arbitro_0:clock
	wire         nios2_custom_instruction_master_multi_slave_translator1_ci_master_clk_en; // nios2_custom_instruction_master_multi_slave_translator1:ci_master_clken -> arbitro_0:clock_en
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator1_ci_master_dataa;  // nios2_custom_instruction_master_multi_slave_translator1:ci_master_dataa -> arbitro_0:dataA
	wire         nios2_custom_instruction_master_multi_slave_translator1_ci_master_reset;  // nios2_custom_instruction_master_multi_slave_translator1:ci_master_reset -> arbitro_0:reset
	wire         nios2_custom_instruction_master_multi_slave_translator1_ci_master_done;   // arbitro_0:done -> nios2_custom_instruction_master_multi_slave_translator1:ci_master_done
	wire  [31:0] nios2_data_master_readdata;                                               // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_waitrequest;                                            // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                                            // nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire  [16:0] nios2_data_master_address;                                                // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                                             // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         nios2_data_master_read;                                                   // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire         nios2_data_master_write;                                                  // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                                              // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                                        // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                                     // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [16:0] nios2_instruction_master_address;                                         // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                                            // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;                      // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;                        // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;                     // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;                         // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;                            // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;                           // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;                       // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;                    // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;                     // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;                         // nios2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;                      // nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;                      // mm_interconnect_0:nios2_debug_mem_slave_debugaccess -> nios2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;                          // mm_interconnect_0:nios2_debug_mem_slave_address -> nios2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;                             // mm_interconnect_0:nios2_debug_mem_slave_read -> nios2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;                       // mm_interconnect_0:nios2_debug_mem_slave_byteenable -> nios2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;                            // mm_interconnect_0:nios2_debug_mem_slave_write -> nios2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;                        // mm_interconnect_0:nios2_debug_mem_slave_writedata -> nios2:debug_mem_slave_writedata
	wire         mm_interconnect_0_memory_s1_chipselect;                                   // mm_interconnect_0:memory_s1_chipselect -> memory:chipselect
	wire  [31:0] mm_interconnect_0_memory_s1_readdata;                                     // memory:readdata -> mm_interconnect_0:memory_s1_readdata
	wire  [12:0] mm_interconnect_0_memory_s1_address;                                      // mm_interconnect_0:memory_s1_address -> memory:address
	wire   [3:0] mm_interconnect_0_memory_s1_byteenable;                                   // mm_interconnect_0:memory_s1_byteenable -> memory:byteenable
	wire         mm_interconnect_0_memory_s1_write;                                        // mm_interconnect_0:memory_s1_write -> memory:write
	wire  [31:0] mm_interconnect_0_memory_s1_writedata;                                    // mm_interconnect_0:memory_s1_writedata -> memory:writedata
	wire         mm_interconnect_0_memory_s1_clken;                                        // mm_interconnect_0:memory_s1_clken -> memory:clken
	wire  [31:0] mm_interconnect_0_pushbutton_s1_readdata;                                 // pushButton:readdata -> mm_interconnect_0:pushButton_s1_readdata
	wire   [1:0] mm_interconnect_0_pushbutton_s1_address;                                  // mm_interconnect_0:pushButton_s1_address -> pushButton:address
	wire         mm_interconnect_0_leds_s1_chipselect;                                     // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                                       // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                                        // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_write;                                          // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                                      // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire         mm_interconnect_0_uart_0_s1_chipselect;                                   // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                                     // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                                      // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;                                         // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                                // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;                                        // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                                    // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire         irq_mapper_receiver0_irq;                                                 // jtag:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                 // uart_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_irq_irq;                                                            // irq_mapper:sender_irq -> nios2:irq
	wire         rst_controller_reset_out_reset;                                           // rst_controller:reset_out -> [irq_mapper:reset, jtag:rst_n, leds:reset_n, memory:reset, mm_interconnect_0:nios2_reset_reset_bridge_in_reset_reset, nios2:reset_n, pushButton:reset_n, rst_translator:in_reset, sysid_qsys_0:reset_n, uart_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                                       // rst_controller:reset_req -> [memory:reset_req, nios2:reset_req, rst_translator:reset_req_in]

	lcd lcd_0 (
		.dataa   (nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // nios_custom_instruction_slave_2.dataa
		.datab   (nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //                                .datab
		.clk     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //                                .clk
		.clk_en  (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //                                .clk_en
		.display (lcd_0_conduit_end_1_readdata),                                             //                   conduit_end_1.readdata
		.rw      (lcd_0_conduit_end_2_writeresponsevalid_n),                                 //                   conduit_end_2.writeresponsevalid_n
		.rs      (lcd_0_conduit_end_3_writeresponsevalid_n),                                 //                   conduit_end_3.writeresponsevalid_n
		.en      (lcd_0_conduit_end_4_writeresponsevalid_n)                                  //                   conduit_end_4.writeresponsevalid_n
	);

	arbitro #(
		.IDLE              (4'b0000),
		.REQUEST           (4'b0001),
		.ANSWER_TIME       (4'b0010),
		.TIMEOUT           (4'b0011),
		.CHECKSUM          (4'b0100),
		.SEND_BACK         (4'b0101),
		.TRYALARM          (5'b00110),
		.c_CLOCK_PERIOD_NS (100)
	) arbitro_0 (
		.clock    (nios2_custom_instruction_master_multi_slave_translator1_ci_master_clk),    // nios_custom_instruction_slave.clk
		.reset    (nios2_custom_instruction_master_multi_slave_translator1_ci_master_reset),  //                              .reset
		.clock_en (nios2_custom_instruction_master_multi_slave_translator1_ci_master_clk_en), //                              .clk_en
		.dataA    (nios2_custom_instruction_master_multi_slave_translator1_ci_master_dataa),  //                              .dataa
		.done     (nios2_custom_instruction_master_multi_slave_translator1_ci_master_done),   //                              .done
		.result   (nios2_custom_instruction_master_multi_slave_translator1_ci_master_result), //                              .result
		.tx       (arbitrotx_writeresponsevalid_n)                                            //                            tx.writeresponsevalid_n
	);

	nios_jtag jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	nios_leds leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_external_connection_export)       // external_connection.export
	);

	nios_memory memory (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),     //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	nios_nios2 nios2 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.E_ci_multi_done                     (nios2_custom_instruction_master_done),                // custom_instruction_master.done
		.E_ci_multi_clk_en                   (nios2_custom_instruction_master_clk_en),              //                          .clk_en
		.E_ci_multi_start                    (nios2_custom_instruction_master_start),               //                          .start
		.E_ci_result                         (nios2_custom_instruction_master_result),              //                          .result
		.D_ci_a                              (nios2_custom_instruction_master_a),                   //                          .a
		.D_ci_b                              (nios2_custom_instruction_master_b),                   //                          .b
		.D_ci_c                              (nios2_custom_instruction_master_c),                   //                          .c
		.D_ci_n                              (nios2_custom_instruction_master_n),                   //                          .n
		.D_ci_readra                         (nios2_custom_instruction_master_readra),              //                          .readra
		.D_ci_readrb                         (nios2_custom_instruction_master_readrb),              //                          .readrb
		.D_ci_writerc                        (nios2_custom_instruction_master_writerc),             //                          .writerc
		.E_ci_dataa                          (nios2_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_datab                          (nios2_custom_instruction_master_datab),               //                          .datab
		.E_ci_multi_clock                    (nios2_custom_instruction_master_clk),                 //                          .clk
		.E_ci_multi_reset                    (nios2_custom_instruction_master_reset),               //                          .reset
		.E_ci_multi_reset_req                (nios2_custom_instruction_master_reset_req),           //                          .reset_req
		.W_ci_estatus                        (nios2_custom_instruction_master_estatus),             //                          .estatus
		.W_ci_ipending                       (nios2_custom_instruction_master_ipending)             //                          .ipending
	);

	nios_pushButton pushbutton (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_pushbutton_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pushbutton_s1_readdata), //                    .readdata
		.in_port  (pushbutton_external_connection_export)     // external_connection.export
	);

	nios_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	nios_uart_0 uart_0 (
		.clk           (clk_clk),                                   //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.rxd           (uart_0_external_connection_rxd),            // external_connection.export
		.txd           (uart_0_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver1_irq)                   //                 irq.irq
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) nios2_custom_instruction_master_translator (
		.ci_slave_dataa            (nios2_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (nios2_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (nios2_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (nios2_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (nios2_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (nios2_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (nios2_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (nios2_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (nios2_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (nios2_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (nios2_custom_instruction_master_ipending),                             //                .ipending
		.ci_slave_estatus          (nios2_custom_instruction_master_estatus),                              //                .estatus
		.ci_slave_multi_clk        (nios2_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_custom_instruction_master_done),                                 //                .done
		.comb_ci_master_dataa      (),                                                                     //  comb_ci_master.dataa
		.comb_ci_master_datab      (),                                                                     //                .datab
		.comb_ci_master_result     (),                                                                     //                .result
		.comb_ci_master_n          (),                                                                     //                .n
		.comb_ci_master_readra     (),                                                                     //                .readra
		.comb_ci_master_readrb     (),                                                                     //                .readrb
		.comb_ci_master_writerc    (),                                                                     //                .writerc
		.comb_ci_master_a          (),                                                                     //                .a
		.comb_ci_master_b          (),                                                                     //                .b
		.comb_ci_master_c          (),                                                                     //                .c
		.comb_ci_master_ipending   (),                                                                     //                .ipending
		.comb_ci_master_estatus    (),                                                                     //                .estatus
		.multi_ci_master_clk       (nios2_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                 //     (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                 //     (terminated)
		.ci_slave_multi_result     (),                                                                     //     (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                          //     (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                 //     (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                 //     (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                 //     (terminated)
		.ci_slave_multi_a          (5'b00000),                                                             //     (terminated)
		.ci_slave_multi_b          (5'b00000),                                                             //     (terminated)
		.ci_slave_multi_c          (5'b00000)                                                              //     (terminated)
	);

	nios_nios2_custom_instruction_master_multi_xconnect nios2_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                     //           .ipending
		.ci_slave_estatus     (),                                                                     //           .estatus
		.ci_slave_clk         (nios2_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_custom_instruction_master_multi_xconnect_ci_master0_done),       //           .done
		.ci_master1_dataa     (nios2_custom_instruction_master_multi_xconnect_ci_master1_dataa),      // ci_master1.dataa
		.ci_master1_datab     (nios2_custom_instruction_master_multi_xconnect_ci_master1_datab),      //           .datab
		.ci_master1_result    (nios2_custom_instruction_master_multi_xconnect_ci_master1_result),     //           .result
		.ci_master1_n         (nios2_custom_instruction_master_multi_xconnect_ci_master1_n),          //           .n
		.ci_master1_readra    (nios2_custom_instruction_master_multi_xconnect_ci_master1_readra),     //           .readra
		.ci_master1_readrb    (nios2_custom_instruction_master_multi_xconnect_ci_master1_readrb),     //           .readrb
		.ci_master1_writerc   (nios2_custom_instruction_master_multi_xconnect_ci_master1_writerc),    //           .writerc
		.ci_master1_a         (nios2_custom_instruction_master_multi_xconnect_ci_master1_a),          //           .a
		.ci_master1_b         (nios2_custom_instruction_master_multi_xconnect_ci_master1_b),          //           .b
		.ci_master1_c         (nios2_custom_instruction_master_multi_xconnect_ci_master1_c),          //           .c
		.ci_master1_ipending  (nios2_custom_instruction_master_multi_xconnect_ci_master1_ipending),   //           .ipending
		.ci_master1_estatus   (nios2_custom_instruction_master_multi_xconnect_ci_master1_estatus),    //           .estatus
		.ci_master1_clk       (nios2_custom_instruction_master_multi_xconnect_ci_master1_clk),        //           .clk
		.ci_master1_reset     (nios2_custom_instruction_master_multi_xconnect_ci_master1_reset),      //           .reset
		.ci_master1_clken     (nios2_custom_instruction_master_multi_xconnect_ci_master1_clk_en),     //           .clk_en
		.ci_master1_reset_req (nios2_custom_instruction_master_multi_xconnect_ci_master1_reset_req),  //           .reset_req
		.ci_master1_start     (nios2_custom_instruction_master_multi_xconnect_ci_master1_start),      //           .start
		.ci_master1_done      (nios2_custom_instruction_master_multi_xconnect_ci_master1_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) nios2_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios2_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios2_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (),                                                                         //          .result
		.ci_master_clk       (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (),                                                                         //          .reset
		.ci_master_n         (),                                                                         // (terminated)
		.ci_master_readra    (),                                                                         // (terminated)
		.ci_master_readrb    (),                                                                         // (terminated)
		.ci_master_writerc   (),                                                                         // (terminated)
		.ci_master_a         (),                                                                         // (terminated)
		.ci_master_b         (),                                                                         // (terminated)
		.ci_master_c         (),                                                                         // (terminated)
		.ci_master_ipending  (),                                                                         // (terminated)
		.ci_master_estatus   (),                                                                         // (terminated)
		.ci_master_reset_req (),                                                                         // (terminated)
		.ci_master_start     (),                                                                         // (terminated)
		.ci_master_done      (1'b0)                                                                      // (terminated)
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios2_custom_instruction_master_multi_slave_translator1 (
		.ci_slave_dataa      (nios2_custom_instruction_master_multi_xconnect_ci_master1_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_custom_instruction_master_multi_xconnect_ci_master1_datab),          //          .datab
		.ci_slave_result     (nios2_custom_instruction_master_multi_xconnect_ci_master1_result),         //          .result
		.ci_slave_n          (nios2_custom_instruction_master_multi_xconnect_ci_master1_n),              //          .n
		.ci_slave_readra     (nios2_custom_instruction_master_multi_xconnect_ci_master1_readra),         //          .readra
		.ci_slave_readrb     (nios2_custom_instruction_master_multi_xconnect_ci_master1_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_custom_instruction_master_multi_xconnect_ci_master1_writerc),        //          .writerc
		.ci_slave_a          (nios2_custom_instruction_master_multi_xconnect_ci_master1_a),              //          .a
		.ci_slave_b          (nios2_custom_instruction_master_multi_xconnect_ci_master1_b),              //          .b
		.ci_slave_c          (nios2_custom_instruction_master_multi_xconnect_ci_master1_c),              //          .c
		.ci_slave_ipending   (nios2_custom_instruction_master_multi_xconnect_ci_master1_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_custom_instruction_master_multi_xconnect_ci_master1_estatus),        //          .estatus
		.ci_slave_clk        (nios2_custom_instruction_master_multi_xconnect_ci_master1_clk),            //          .clk
		.ci_slave_clken      (nios2_custom_instruction_master_multi_xconnect_ci_master1_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_custom_instruction_master_multi_xconnect_ci_master1_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_custom_instruction_master_multi_xconnect_ci_master1_reset),          //          .reset
		.ci_slave_start      (nios2_custom_instruction_master_multi_xconnect_ci_master1_start),          //          .start
		.ci_slave_done       (nios2_custom_instruction_master_multi_xconnect_ci_master1_done),           //          .done
		.ci_master_dataa     (nios2_custom_instruction_master_multi_slave_translator1_ci_master_dataa),  // ci_master.dataa
		.ci_master_result    (nios2_custom_instruction_master_multi_slave_translator1_ci_master_result), //          .result
		.ci_master_clk       (nios2_custom_instruction_master_multi_slave_translator1_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_custom_instruction_master_multi_slave_translator1_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_custom_instruction_master_multi_slave_translator1_ci_master_reset),  //          .reset
		.ci_master_done      (nios2_custom_instruction_master_multi_slave_translator1_ci_master_done),   //          .done
		.ci_master_datab     (),                                                                         // (terminated)
		.ci_master_n         (),                                                                         // (terminated)
		.ci_master_readra    (),                                                                         // (terminated)
		.ci_master_readrb    (),                                                                         // (terminated)
		.ci_master_writerc   (),                                                                         // (terminated)
		.ci_master_a         (),                                                                         // (terminated)
		.ci_master_b         (),                                                                         // (terminated)
		.ci_master_c         (),                                                                         // (terminated)
		.ci_master_ipending  (),                                                                         // (terminated)
		.ci_master_estatus   (),                                                                         // (terminated)
		.ci_master_reset_req (),                                                                         // (terminated)
		.ci_master_start     ()                                                                          // (terminated)
	);

	nios_mm_interconnect_0 mm_interconnect_0 (
		.Clk_clk_clk                             (clk_clk),                                               //                           Clk_clk.clk
		.nios2_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // nios2_reset_reset_bridge_in_reset.reset
		.nios2_data_master_address               (nios2_data_master_address),                             //                 nios2_data_master.address
		.nios2_data_master_waitrequest           (nios2_data_master_waitrequest),                         //                                  .waitrequest
		.nios2_data_master_byteenable            (nios2_data_master_byteenable),                          //                                  .byteenable
		.nios2_data_master_read                  (nios2_data_master_read),                                //                                  .read
		.nios2_data_master_readdata              (nios2_data_master_readdata),                            //                                  .readdata
		.nios2_data_master_write                 (nios2_data_master_write),                               //                                  .write
		.nios2_data_master_writedata             (nios2_data_master_writedata),                           //                                  .writedata
		.nios2_data_master_debugaccess           (nios2_data_master_debugaccess),                         //                                  .debugaccess
		.nios2_instruction_master_address        (nios2_instruction_master_address),                      //          nios2_instruction_master.address
		.nios2_instruction_master_waitrequest    (nios2_instruction_master_waitrequest),                  //                                  .waitrequest
		.nios2_instruction_master_read           (nios2_instruction_master_read),                         //                                  .read
		.nios2_instruction_master_readdata       (nios2_instruction_master_readdata),                     //                                  .readdata
		.jtag_avalon_jtag_slave_address          (mm_interconnect_0_jtag_avalon_jtag_slave_address),      //            jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write            (mm_interconnect_0_jtag_avalon_jtag_slave_write),        //                                  .write
		.jtag_avalon_jtag_slave_read             (mm_interconnect_0_jtag_avalon_jtag_slave_read),         //                                  .read
		.jtag_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),     //                                  .readdata
		.jtag_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),    //                                  .writedata
		.jtag_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),  //                                  .waitrequest
		.jtag_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),   //                                  .chipselect
		.leds_s1_address                         (mm_interconnect_0_leds_s1_address),                     //                           leds_s1.address
		.leds_s1_write                           (mm_interconnect_0_leds_s1_write),                       //                                  .write
		.leds_s1_readdata                        (mm_interconnect_0_leds_s1_readdata),                    //                                  .readdata
		.leds_s1_writedata                       (mm_interconnect_0_leds_s1_writedata),                   //                                  .writedata
		.leds_s1_chipselect                      (mm_interconnect_0_leds_s1_chipselect),                  //                                  .chipselect
		.memory_s1_address                       (mm_interconnect_0_memory_s1_address),                   //                         memory_s1.address
		.memory_s1_write                         (mm_interconnect_0_memory_s1_write),                     //                                  .write
		.memory_s1_readdata                      (mm_interconnect_0_memory_s1_readdata),                  //                                  .readdata
		.memory_s1_writedata                     (mm_interconnect_0_memory_s1_writedata),                 //                                  .writedata
		.memory_s1_byteenable                    (mm_interconnect_0_memory_s1_byteenable),                //                                  .byteenable
		.memory_s1_chipselect                    (mm_interconnect_0_memory_s1_chipselect),                //                                  .chipselect
		.memory_s1_clken                         (mm_interconnect_0_memory_s1_clken),                     //                                  .clken
		.nios2_debug_mem_slave_address           (mm_interconnect_0_nios2_debug_mem_slave_address),       //             nios2_debug_mem_slave.address
		.nios2_debug_mem_slave_write             (mm_interconnect_0_nios2_debug_mem_slave_write),         //                                  .write
		.nios2_debug_mem_slave_read              (mm_interconnect_0_nios2_debug_mem_slave_read),          //                                  .read
		.nios2_debug_mem_slave_readdata          (mm_interconnect_0_nios2_debug_mem_slave_readdata),      //                                  .readdata
		.nios2_debug_mem_slave_writedata         (mm_interconnect_0_nios2_debug_mem_slave_writedata),     //                                  .writedata
		.nios2_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_debug_mem_slave_byteenable),    //                                  .byteenable
		.nios2_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),   //                                  .waitrequest
		.nios2_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),   //                                  .debugaccess
		.pushButton_s1_address                   (mm_interconnect_0_pushbutton_s1_address),               //                     pushButton_s1.address
		.pushButton_s1_readdata                  (mm_interconnect_0_pushbutton_s1_readdata),              //                                  .readdata
		.sysid_qsys_0_control_slave_address      (mm_interconnect_0_sysid_qsys_0_control_slave_address),  //        sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata     (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), //                                  .readdata
		.uart_0_s1_address                       (mm_interconnect_0_uart_0_s1_address),                   //                         uart_0_s1.address
		.uart_0_s1_write                         (mm_interconnect_0_uart_0_s1_write),                     //                                  .write
		.uart_0_s1_read                          (mm_interconnect_0_uart_0_s1_read),                      //                                  .read
		.uart_0_s1_readdata                      (mm_interconnect_0_uart_0_s1_readdata),                  //                                  .readdata
		.uart_0_s1_writedata                     (mm_interconnect_0_uart_0_s1_writedata),                 //                                  .writedata
		.uart_0_s1_begintransfer                 (mm_interconnect_0_uart_0_s1_begintransfer),             //                                  .begintransfer
		.uart_0_s1_chipselect                    (mm_interconnect_0_uart_0_s1_chipselect)                 //                                  .chipselect
	);

	nios_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_debug_reset_request_reset),    // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
